configuration of vectorgate_struc_cfg of vectorgate is

	for struc
		end for;
	end vectorgate_struc_cfg;
