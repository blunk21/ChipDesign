library IEEE;
use IEEE.std_logic_1164.all;

entity tb_decoder is
end tb_decoder;