configuration tb_xorgate_sim_cfg of tb_xorgate is
	for sim
	end for;
end tb_xorgate_sim_cfg;
