library IEEE;
use IEEE.std_logic_1164.all;

entity tb_xorgate is
end tb_xorgate;
