library IEEE;
use IEEE.std_logic_1164.all;



entity xorgate is
	port (a_i : in std_logic;
	      b_i : in std_logic;
    	      xor_o : out std_logic);
end xorgate;	






